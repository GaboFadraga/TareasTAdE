
Started : "Check Syntax for counter".
Running xst...
Command Line: xst -intstyle ise -ifn {/home/ise/Gabriel/Desktop/Tareas TAdE/Pregunta1Preparacion/counter.xst} -ofn counter.stx

=========================================================================
*                          HDL Compilation                              *
=========================================================================
Compiling vhdl file "/home/ise/Gabriel/Desktop/Tareas TAdE/Pregunta1Preparacion/ej1.vhd" in Library work.
Architecture behavioral of Entity counter is up to date.

Process "Check Syntax" completed successfully
